module top_1598227639_809568180_776209382_1234615 (n1, n2, n4, n5, n7);
  input n1, n2, n4, n5;
  output n7;
  xnor_6 g0(n1,n2,n3);
  xnor_6 g1(n4,n5,n6);
  xnor_6 g2(n3,n6,n7);
endmodule
