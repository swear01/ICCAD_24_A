module top_809960632_810038711_1598227639_893650103(n1, n2, n3);
  input n1, n2;
  output n3;
  and_1 g0 ( n1 , n2 , n3 ) ;
endmodule
