module top_1598227639_809568180_776209382_1234615 (n2, n4, n12, n18, n22, n34, n35, n51, n57, n67, n72, n75, n78, n80, n6, n9, n42, n48, n56, n65, n68, n77);
  input n2, n4, n12, n18, n22, n34, n35, n51, n57, n67, n72, n75, n78, n80;
  output n6, n9, n42, n48, n56, n65, n68, n77;
  or_4 g0(n86,n73,n77);
  xnor_5 g1(n45,n53,n5);
  xor_4 g2(n61,n30,n9);
  nor_3 g3(n12,n27,n40);
  not_11 g4(n10,n16);
  not_4 g5(n84,n81);
  and_1 g6(n34,n44,n31);
  or_1 g7(n80,n2,n26);
  and_3 g8(n72,n67,n58);
  not_4 g9(n2,n24);
  or_4 g10(n21,n78,n14);
  and_7 g11(n39,n1,n79);
  or_3 g12(n80,n67,n20);
  nor_8 g13(n84,n76,n7);
  and_5 g14(n72,n57,n52);
  and_3 g15(n28,n36,n50);
  not_5 g16(n45,n15);
  xnor_1 g17(n0,n50,n69);
  nand_2 g18(n72,n4,n3);
  and_8 g19(n22,n20,n43);
  and_6 g20(n53,n16,n27);
  not_13 g21(n4,n21);
  or_3 g22(n37,n12,n60);
  and_7 g23(n55,n70,n1);
  not_11 g24(n67,n88);
  and_6 g25(n18,n26,n87);
  not_4 g26(n63,n48);
  not_13 g27(n57,n71);
  xnor_4 g28(n60,n5,n6);
  nor_6 g29(n37,n77,n33);
  and_6 g30(n35,n25,n59);
  and_2 g31(n54,n43,n45);
  or_1 g32(n52,n64,n55);
  not_9 g33(n75,n29);
  nor_2 g34(n29,n4,n74);
  or_1 g35(n90,n11,n86);
  or_2 g36(n66,n45,n73);
  xor_1 g37(n40,n69,n42);
  xor_2 g38(n19,n82,n65);
  and_3 g39(n9,n65,n89);
  not_5 g40(n51,n37);
  and_2 g41(n14,n59,n90);
  or_1 g42(n80,n4,n25);
  and_2 g43(n3,n38,n49);
  and_8 g44(n51,n15,n10);
  nor_7 g45(n12,n7,n61);
  or_3 g46(n33,n63,n68);
  or_2 g47(n11,n47,n70);
  nor_2 g48(n18,n23,n36);
  or_1 g49(n71,n78,n46);
  nor_8 g50(n90,n1,n32);
  or_2 g51(n11,n81,n39);
  nor_7 g52(n29,n57,n13);
  xor_2 g53(n90,n49,n82);
  and_4 g54(n8,n89,n56);
  xnor_1 g55(n11,n55,n30);
  or_4 g56(n22,n83,n41);
  or_4 g57(n88,n78,n54);
  not_3 g58(n72,n17);
  nor_8 g59(n12,n79,n19);
  nor_6 g60(n35,n74,n38);
  and_7 g61(n46,n31,n11);
  nor_1 g62(n29,n2,n23);
  or_7 g63(n80,n57,n44);
  or_1 g64(n50,n62,n76);
  and_6 g65(n85,n87,n66);
  or_4 g66(n58,n41,n53);
  or_7 g67(n24,n78,n85);
  nor_2 g68(n29,n67,n83);
  not_12 g69(n66,n0);
  not_10 g70(n76,n47);
  or_3 g71(n49,n32,n63);
  nor_5 g72(n53,n66,n62);
  and_6 g73(n6,n42,n8);
  and_6 g74(n0,n10,n84);
  or_5 g75(n34,n13,n64);
  or_1 g76(n17,n24,n28);
endmodule
