module top_809960632_810038711_1598227639_893650103 (n1,n2,n3);
  input n1_1,n2,n4,n5;
  output n7;
  or_8 g0(n1_1,n2,n3);
  or_8 g1(n4,n5,n6);
  or_8 g2(n3,n6,n7);
endmodule